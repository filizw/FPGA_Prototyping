`timescale 1ns / 1ps

// 12-to-4 priority encoder
module prio_enc(
    input [11:0] r,
    output reg [3:0] y
    );

	always @*
	begin
		casez(r)
			12'b1???????????: y = 4'd12;
			12'b01??????????: y = 4'd11;
			12'b001?????????: y = 4'd10;
			12'b0001????????: y = 4'd9;
			12'b00001???????: y = 4'd8;
			12'b000001??????: y = 4'd7;
			12'b0000001?????: y = 4'd6;
			12'b00000001????: y = 4'd5;
			12'b000000001???: y = 4'd4;
			12'b0000000001??: y = 4'd3;
			12'b00000000001?: y = 4'd2;
			12'b000000000001: y = 4'd1;
			default: y = 4'd0;
		endcase
	end

endmodule
